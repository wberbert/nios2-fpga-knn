// nios2_sopc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios2_sopc (
		input  wire        clk50_0_clk,                             //                          clk50_0.clk
		input  wire [15:0] knn_classe_prevista_distancia_in_export, // knn_classe_prevista_distancia_in.export
		input  wire [15:0] knn_classe_prevista_in_export,           //           knn_classe_prevista_in.export
		input  wire        knn_classe_prevista_pronto_in_export,    //    knn_classe_prevista_pronto_in.export
		output wire [7:0]  knn_dados_atributo_out_export,           //           knn_dados_atributo_out.export
		output wire        knn_dados_pronto_out_export,             //             knn_dados_pronto_out.export
		output wire [15:0] knn_dados_valor_out_export,              //              knn_dados_valor_out.export
		output wire [3:0]  knn_k_out_export,                        //                        knn_k_out.export
		output wire        knn_reset_out_export,                    //                    knn_reset_out.export
		output wire        knn_treinamento_out_export,              //              knn_treinamento_out.export
		output wire [7:0]  pio_0_external_connection_export,        //        pio_0_external_connection.export
		input  wire        reset_clk50_0_reset_n,                   //                    reset_clk50_0.reset_n
		input  wire        rs232_0_external_interface_RXD,          //       rs232_0_external_interface.RXD
		output wire        rs232_0_external_interface_TXD,          //                                 .TXD
		output wire [12:0] sdram_0_wire_addr,                       //                     sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                         //                                 .ba
		output wire        sdram_0_wire_cas_n,                      //                                 .cas_n
		output wire        sdram_0_wire_cke,                        //                                 .cke
		output wire        sdram_0_wire_cs_n,                       //                                 .cs_n
		inout  wire [31:0] sdram_0_wire_dq,                         //                                 .dq
		output wire [3:0]  sdram_0_wire_dqm,                        //                                 .dqm
		output wire        sdram_0_wire_ras_n,                      //                                 .ras_n
		output wire        sdram_0_wire_we_n,                       //                                 .we_n
		input  wire        usb_0_external_interface_INT1,           //         usb_0_external_interface.INT1
		inout  wire [15:0] usb_0_external_interface_DATA,           //                                 .DATA
		output wire        usb_0_external_interface_RST_N,          //                                 .RST_N
		output wire [1:0]  usb_0_external_interface_ADDR,           //                                 .ADDR
		output wire        usb_0_external_interface_CS_N,           //                                 .CS_N
		output wire        usb_0_external_interface_RD_N,           //                                 .RD_N
		output wire        usb_0_external_interface_WR_N,           //                                 .WR_N
		input  wire        usb_0_external_interface_INT0,           //                                 .INT0
		output wire        vga_0_external_interface_CLK,            //         vga_0_external_interface.CLK
		output wire        vga_0_external_interface_HS,             //                                 .HS
		output wire        vga_0_external_interface_VS,             //                                 .VS
		output wire        vga_0_external_interface_BLANK,          //                                 .BLANK
		output wire        vga_0_external_interface_SYNC,           //                                 .SYNC
		output wire [7:0]  vga_0_external_interface_R,              //                                 .R
		output wire [7:0]  vga_0_external_interface_G,              //                                 .G
		output wire [7:0]  vga_0_external_interface_B               //                                 .B
	);

	wire         vga_buffer_0_avalon_char_source_valid;                               // VGA_BUFFER_0:stream_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire  [29:0] vga_buffer_0_avalon_char_source_data;                                // VGA_BUFFER_0:stream_data -> video_dual_clock_buffer_0:stream_in_data
	wire         vga_buffer_0_avalon_char_source_ready;                               // video_dual_clock_buffer_0:stream_in_ready -> VGA_BUFFER_0:stream_ready
	wire         vga_buffer_0_avalon_char_source_startofpacket;                       // VGA_BUFFER_0:stream_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire         vga_buffer_0_avalon_char_source_endofpacket;                         // VGA_BUFFER_0:stream_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;             // video_dual_clock_buffer_0:stream_out_valid -> VGA_0:valid
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;              // video_dual_clock_buffer_0:stream_out_data -> VGA_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;             // VGA_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;     // video_dual_clock_buffer_0:stream_out_startofpacket -> VGA_0:startofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;       // video_dual_clock_buffer_0:stream_out_endofpacket -> VGA_0:endofpacket
	wire         vga_pll_0_c0_clk;                                                    // VGA_PLL_0:c0 -> [VGA_0:clk, VGA_BUFFER_0:clk, mm_interconnect_0:VGA_PLL_0_c0_clk, rst_controller_001:clk, rst_controller_002:clk, video_dual_clock_buffer_0:clk_stream_in, video_dual_clock_buffer_0:clk_stream_out]
	wire  [31:0] nios2_0_data_master_readdata;                                        // mm_interconnect_0:NIOS2_0_data_master_readdata -> NIOS2_0:d_readdata
	wire         nios2_0_data_master_waitrequest;                                     // mm_interconnect_0:NIOS2_0_data_master_waitrequest -> NIOS2_0:d_waitrequest
	wire         nios2_0_data_master_debugaccess;                                     // NIOS2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_0_data_master_debugaccess
	wire  [27:0] nios2_0_data_master_address;                                         // NIOS2_0:d_address -> mm_interconnect_0:NIOS2_0_data_master_address
	wire   [3:0] nios2_0_data_master_byteenable;                                      // NIOS2_0:d_byteenable -> mm_interconnect_0:NIOS2_0_data_master_byteenable
	wire         nios2_0_data_master_read;                                            // NIOS2_0:d_read -> mm_interconnect_0:NIOS2_0_data_master_read
	wire         nios2_0_data_master_readdatavalid;                                   // mm_interconnect_0:NIOS2_0_data_master_readdatavalid -> NIOS2_0:d_readdatavalid
	wire         nios2_0_data_master_write;                                           // NIOS2_0:d_write -> mm_interconnect_0:NIOS2_0_data_master_write
	wire  [31:0] nios2_0_data_master_writedata;                                       // NIOS2_0:d_writedata -> mm_interconnect_0:NIOS2_0_data_master_writedata
	wire  [31:0] nios2_0_instruction_master_readdata;                                 // mm_interconnect_0:NIOS2_0_instruction_master_readdata -> NIOS2_0:i_readdata
	wire         nios2_0_instruction_master_waitrequest;                              // mm_interconnect_0:NIOS2_0_instruction_master_waitrequest -> NIOS2_0:i_waitrequest
	wire  [27:0] nios2_0_instruction_master_address;                                  // NIOS2_0:i_address -> mm_interconnect_0:NIOS2_0_instruction_master_address
	wire         nios2_0_instruction_master_read;                                     // NIOS2_0:i_read -> mm_interconnect_0:NIOS2_0_instruction_master_read
	wire         nios2_0_instruction_master_readdatavalid;                            // mm_interconnect_0:NIOS2_0_instruction_master_readdatavalid -> NIOS2_0:i_readdatavalid
	wire         mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_chipselect -> VGA_BUFFER_0:buf_chipselect
	wire   [7:0] mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_readdata;    // VGA_BUFFER_0:buf_readdata -> mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_waitrequest; // VGA_BUFFER_0:buf_waitrequest -> mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_address;     // mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_address -> VGA_BUFFER_0:buf_address
	wire         mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_read;        // mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_read -> VGA_BUFFER_0:buf_read
	wire   [0:0] mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_byteenable -> VGA_BUFFER_0:buf_byteenable
	wire         mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_write;       // mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_write -> VGA_BUFFER_0:buf_write
	wire   [7:0] mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:VGA_BUFFER_0_avalon_char_buffer_slave_writedata -> VGA_BUFFER_0:buf_writedata
	wire         mm_interconnect_0_jtag_0_avalon_jtag_slave_chipselect;               // mm_interconnect_0:JTAG_0_avalon_jtag_slave_chipselect -> JTAG_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_0_avalon_jtag_slave_readdata;                 // JTAG_0:av_readdata -> mm_interconnect_0:JTAG_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_0_avalon_jtag_slave_waitrequest;              // JTAG_0:av_waitrequest -> mm_interconnect_0:JTAG_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_0_avalon_jtag_slave_address;                  // mm_interconnect_0:JTAG_0_avalon_jtag_slave_address -> JTAG_0:av_address
	wire         mm_interconnect_0_jtag_0_avalon_jtag_slave_read;                     // mm_interconnect_0:JTAG_0_avalon_jtag_slave_read -> JTAG_0:av_read_n
	wire         mm_interconnect_0_jtag_0_avalon_jtag_slave_write;                    // mm_interconnect_0:JTAG_0_avalon_jtag_slave_write -> JTAG_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_0_avalon_jtag_slave_writedata;                // mm_interconnect_0:JTAG_0_avalon_jtag_slave_writedata -> JTAG_0:av_writedata
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect;             // mm_interconnect_0:RS232_0_avalon_rs232_slave_chipselect -> RS232_0:chipselect
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata;               // RS232_0:readdata -> mm_interconnect_0:RS232_0_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_address;                // mm_interconnect_0:RS232_0_avalon_rs232_slave_address -> RS232_0:address
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_read;                   // mm_interconnect_0:RS232_0_avalon_rs232_slave_read -> RS232_0:read
	wire   [3:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable;             // mm_interconnect_0:RS232_0_avalon_rs232_slave_byteenable -> RS232_0:byteenable
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_write;                  // mm_interconnect_0:RS232_0_avalon_rs232_slave_write -> RS232_0:write
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata;              // mm_interconnect_0:RS232_0_avalon_rs232_slave_writedata -> RS232_0:writedata
	wire         mm_interconnect_0_usb_0_avalon_usb_slave_chipselect;                 // mm_interconnect_0:USB_0_avalon_usb_slave_chipselect -> USB_0:chipselect
	wire  [15:0] mm_interconnect_0_usb_0_avalon_usb_slave_readdata;                   // USB_0:readdata -> mm_interconnect_0:USB_0_avalon_usb_slave_readdata
	wire   [1:0] mm_interconnect_0_usb_0_avalon_usb_slave_address;                    // mm_interconnect_0:USB_0_avalon_usb_slave_address -> USB_0:address
	wire         mm_interconnect_0_usb_0_avalon_usb_slave_read;                       // mm_interconnect_0:USB_0_avalon_usb_slave_read -> USB_0:read
	wire         mm_interconnect_0_usb_0_avalon_usb_slave_write;                      // mm_interconnect_0:USB_0_avalon_usb_slave_write -> USB_0:write
	wire  [15:0] mm_interconnect_0_usb_0_avalon_usb_slave_writedata;                  // mm_interconnect_0:USB_0_avalon_usb_slave_writedata -> USB_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_0_debug_mem_slave_readdata;                  // NIOS2_0:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest;               // NIOS2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess;               // mm_interconnect_0:NIOS2_0_debug_mem_slave_debugaccess -> NIOS2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_0_debug_mem_slave_address;                   // mm_interconnect_0:NIOS2_0_debug_mem_slave_address -> NIOS2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_read;                      // mm_interconnect_0:NIOS2_0_debug_mem_slave_read -> NIOS2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_0_debug_mem_slave_byteenable;                // mm_interconnect_0:NIOS2_0_debug_mem_slave_byteenable -> NIOS2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_write;                     // mm_interconnect_0:NIOS2_0_debug_mem_slave_write -> NIOS2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_0_debug_mem_slave_writedata;                 // mm_interconnect_0:NIOS2_0_debug_mem_slave_writedata -> NIOS2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_vga_pll_0_pll_slave_readdata;                      // VGA_PLL_0:readdata -> mm_interconnect_0:VGA_PLL_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_pll_0_pll_slave_address;                       // mm_interconnect_0:VGA_PLL_0_pll_slave_address -> VGA_PLL_0:address
	wire         mm_interconnect_0_vga_pll_0_pll_slave_read;                          // mm_interconnect_0:VGA_PLL_0_pll_slave_read -> VGA_PLL_0:read
	wire         mm_interconnect_0_vga_pll_0_pll_slave_write;                         // mm_interconnect_0:VGA_PLL_0_pll_slave_write -> VGA_PLL_0:write
	wire  [31:0] mm_interconnect_0_vga_pll_0_pll_slave_writedata;                     // mm_interconnect_0:VGA_PLL_0_pll_slave_writedata -> VGA_PLL_0:writedata
	wire         mm_interconnect_0_mmu_0_s1_chipselect;                               // mm_interconnect_0:MMU_0_s1_chipselect -> MMU_0:chipselect
	wire  [31:0] mm_interconnect_0_mmu_0_s1_readdata;                                 // MMU_0:readdata -> mm_interconnect_0:MMU_0_s1_readdata
	wire   [7:0] mm_interconnect_0_mmu_0_s1_address;                                  // mm_interconnect_0:MMU_0_s1_address -> MMU_0:address
	wire   [3:0] mm_interconnect_0_mmu_0_s1_byteenable;                               // mm_interconnect_0:MMU_0_s1_byteenable -> MMU_0:byteenable
	wire         mm_interconnect_0_mmu_0_s1_write;                                    // mm_interconnect_0:MMU_0_s1_write -> MMU_0:write
	wire  [31:0] mm_interconnect_0_mmu_0_s1_writedata;                                // mm_interconnect_0:MMU_0_s1_writedata -> MMU_0:writedata
	wire         mm_interconnect_0_mmu_0_s1_clken;                                    // mm_interconnect_0:MMU_0_s1_clken -> MMU_0:clken
	wire         mm_interconnect_0_sdram_0_s1_chipselect;                             // mm_interconnect_0:SDRAM_0_s1_chipselect -> SDRAM_0:az_cs
	wire  [31:0] mm_interconnect_0_sdram_0_s1_readdata;                               // SDRAM_0:za_data -> mm_interconnect_0:SDRAM_0_s1_readdata
	wire         mm_interconnect_0_sdram_0_s1_waitrequest;                            // SDRAM_0:za_waitrequest -> mm_interconnect_0:SDRAM_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_0_s1_address;                                // mm_interconnect_0:SDRAM_0_s1_address -> SDRAM_0:az_addr
	wire         mm_interconnect_0_sdram_0_s1_read;                                   // mm_interconnect_0:SDRAM_0_s1_read -> SDRAM_0:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_0_s1_byteenable;                             // mm_interconnect_0:SDRAM_0_s1_byteenable -> SDRAM_0:az_be_n
	wire         mm_interconnect_0_sdram_0_s1_readdatavalid;                          // SDRAM_0:za_valid -> mm_interconnect_0:SDRAM_0_s1_readdatavalid
	wire         mm_interconnect_0_sdram_0_s1_write;                                  // mm_interconnect_0:SDRAM_0_s1_write -> SDRAM_0:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_0_s1_writedata;                              // mm_interconnect_0:SDRAM_0_s1_writedata -> SDRAM_0:az_data
	wire         mm_interconnect_0_pio_0_s1_chipselect;                               // mm_interconnect_0:PIO_0_s1_chipselect -> PIO_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                                 // PIO_0:readdata -> mm_interconnect_0:PIO_0_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_0_s1_address;                                  // mm_interconnect_0:PIO_0_s1_address -> PIO_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                                    // mm_interconnect_0:PIO_0_s1_write -> PIO_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                                // mm_interconnect_0:PIO_0_s1_writedata -> PIO_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                             // mm_interconnect_0:TIMER_1_s1_chipselect -> TIMER_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                               // TIMER_1:readdata -> mm_interconnect_0:TIMER_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                                // mm_interconnect_0:TIMER_1_s1_address -> TIMER_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                                  // mm_interconnect_0:TIMER_1_s1_write -> TIMER_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                              // mm_interconnect_0:TIMER_1_s1_writedata -> TIMER_1:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                             // mm_interconnect_0:TIMER_0_s1_chipselect -> TIMER_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                               // TIMER_0:readdata -> mm_interconnect_0:TIMER_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                // mm_interconnect_0:TIMER_0_s1_address -> TIMER_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                  // mm_interconnect_0:TIMER_0_s1_write -> TIMER_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                              // mm_interconnect_0:TIMER_0_s1_writedata -> TIMER_0:writedata
	wire         mm_interconnect_0_po_knn_dados_s1_chipselect;                        // mm_interconnect_0:PO_KNN_DADOS_s1_chipselect -> PO_KNN_DADOS:chipselect
	wire  [31:0] mm_interconnect_0_po_knn_dados_s1_readdata;                          // PO_KNN_DADOS:readdata -> mm_interconnect_0:PO_KNN_DADOS_s1_readdata
	wire   [1:0] mm_interconnect_0_po_knn_dados_s1_address;                           // mm_interconnect_0:PO_KNN_DADOS_s1_address -> PO_KNN_DADOS:address
	wire         mm_interconnect_0_po_knn_dados_s1_write;                             // mm_interconnect_0:PO_KNN_DADOS_s1_write -> PO_KNN_DADOS:write_n
	wire  [31:0] mm_interconnect_0_po_knn_dados_s1_writedata;                         // mm_interconnect_0:PO_KNN_DADOS_s1_writedata -> PO_KNN_DADOS:writedata
	wire         mm_interconnect_0_po_knn_dados_pronto_s1_chipselect;                 // mm_interconnect_0:PO_KNN_DADOS_PRONTO_s1_chipselect -> PO_KNN_DADOS_PRONTO:chipselect
	wire  [31:0] mm_interconnect_0_po_knn_dados_pronto_s1_readdata;                   // PO_KNN_DADOS_PRONTO:readdata -> mm_interconnect_0:PO_KNN_DADOS_PRONTO_s1_readdata
	wire   [1:0] mm_interconnect_0_po_knn_dados_pronto_s1_address;                    // mm_interconnect_0:PO_KNN_DADOS_PRONTO_s1_address -> PO_KNN_DADOS_PRONTO:address
	wire         mm_interconnect_0_po_knn_dados_pronto_s1_write;                      // mm_interconnect_0:PO_KNN_DADOS_PRONTO_s1_write -> PO_KNN_DADOS_PRONTO:write_n
	wire  [31:0] mm_interconnect_0_po_knn_dados_pronto_s1_writedata;                  // mm_interconnect_0:PO_KNN_DADOS_PRONTO_s1_writedata -> PO_KNN_DADOS_PRONTO:writedata
	wire  [31:0] mm_interconnect_0_pi_knn_classe_prevista_s1_readdata;                // PI_KNN_CLASSE_PREVISTA:readdata -> mm_interconnect_0:PI_KNN_CLASSE_PREVISTA_s1_readdata
	wire   [1:0] mm_interconnect_0_pi_knn_classe_prevista_s1_address;                 // mm_interconnect_0:PI_KNN_CLASSE_PREVISTA_s1_address -> PI_KNN_CLASSE_PREVISTA:address
	wire  [31:0] mm_interconnect_0_pi_knn_classe_prevista_pronto_s1_readdata;         // PI_KNN_CLASSE_PREVISTA_PRONTO:readdata -> mm_interconnect_0:PI_KNN_CLASSE_PREVISTA_PRONTO_s1_readdata
	wire   [1:0] mm_interconnect_0_pi_knn_classe_prevista_pronto_s1_address;          // mm_interconnect_0:PI_KNN_CLASSE_PREVISTA_PRONTO_s1_address -> PI_KNN_CLASSE_PREVISTA_PRONTO:address
	wire         mm_interconnect_0_po_knn_dados_atributo_s1_chipselect;               // mm_interconnect_0:PO_KNN_DADOS_ATRIBUTO_s1_chipselect -> PO_KNN_DADOS_ATRIBUTO:chipselect
	wire  [31:0] mm_interconnect_0_po_knn_dados_atributo_s1_readdata;                 // PO_KNN_DADOS_ATRIBUTO:readdata -> mm_interconnect_0:PO_KNN_DADOS_ATRIBUTO_s1_readdata
	wire   [1:0] mm_interconnect_0_po_knn_dados_atributo_s1_address;                  // mm_interconnect_0:PO_KNN_DADOS_ATRIBUTO_s1_address -> PO_KNN_DADOS_ATRIBUTO:address
	wire         mm_interconnect_0_po_knn_dados_atributo_s1_write;                    // mm_interconnect_0:PO_KNN_DADOS_ATRIBUTO_s1_write -> PO_KNN_DADOS_ATRIBUTO:write_n
	wire  [31:0] mm_interconnect_0_po_knn_dados_atributo_s1_writedata;                // mm_interconnect_0:PO_KNN_DADOS_ATRIBUTO_s1_writedata -> PO_KNN_DADOS_ATRIBUTO:writedata
	wire         mm_interconnect_0_po_knn_treinamento_s1_chipselect;                  // mm_interconnect_0:PO_KNN_TREINAMENTO_s1_chipselect -> PO_KNN_TREINAMENTO:chipselect
	wire  [31:0] mm_interconnect_0_po_knn_treinamento_s1_readdata;                    // PO_KNN_TREINAMENTO:readdata -> mm_interconnect_0:PO_KNN_TREINAMENTO_s1_readdata
	wire   [1:0] mm_interconnect_0_po_knn_treinamento_s1_address;                     // mm_interconnect_0:PO_KNN_TREINAMENTO_s1_address -> PO_KNN_TREINAMENTO:address
	wire         mm_interconnect_0_po_knn_treinamento_s1_write;                       // mm_interconnect_0:PO_KNN_TREINAMENTO_s1_write -> PO_KNN_TREINAMENTO:write_n
	wire  [31:0] mm_interconnect_0_po_knn_treinamento_s1_writedata;                   // mm_interconnect_0:PO_KNN_TREINAMENTO_s1_writedata -> PO_KNN_TREINAMENTO:writedata
	wire         mm_interconnect_0_po_knn_reset_s1_chipselect;                        // mm_interconnect_0:PO_KNN_RESET_s1_chipselect -> PO_KNN_RESET:chipselect
	wire  [31:0] mm_interconnect_0_po_knn_reset_s1_readdata;                          // PO_KNN_RESET:readdata -> mm_interconnect_0:PO_KNN_RESET_s1_readdata
	wire   [1:0] mm_interconnect_0_po_knn_reset_s1_address;                           // mm_interconnect_0:PO_KNN_RESET_s1_address -> PO_KNN_RESET:address
	wire         mm_interconnect_0_po_knn_reset_s1_write;                             // mm_interconnect_0:PO_KNN_RESET_s1_write -> PO_KNN_RESET:write_n
	wire  [31:0] mm_interconnect_0_po_knn_reset_s1_writedata;                         // mm_interconnect_0:PO_KNN_RESET_s1_writedata -> PO_KNN_RESET:writedata
	wire         mm_interconnect_0_po_knn_k_s1_chipselect;                            // mm_interconnect_0:PO_KNN_K_s1_chipselect -> PO_KNN_K:chipselect
	wire  [31:0] mm_interconnect_0_po_knn_k_s1_readdata;                              // PO_KNN_K:readdata -> mm_interconnect_0:PO_KNN_K_s1_readdata
	wire   [1:0] mm_interconnect_0_po_knn_k_s1_address;                               // mm_interconnect_0:PO_KNN_K_s1_address -> PO_KNN_K:address
	wire         mm_interconnect_0_po_knn_k_s1_write;                                 // mm_interconnect_0:PO_KNN_K_s1_write -> PO_KNN_K:write_n
	wire  [31:0] mm_interconnect_0_po_knn_k_s1_writedata;                             // mm_interconnect_0:PO_KNN_K_s1_writedata -> PO_KNN_K:writedata
	wire  [31:0] mm_interconnect_0_pi_knn_classe_prevista_distancia_s1_readdata;      // PI_KNN_CLASSE_PREVISTA_DISTANCIA:readdata -> mm_interconnect_0:PI_KNN_CLASSE_PREVISTA_DISTANCIA_s1_readdata
	wire   [1:0] mm_interconnect_0_pi_knn_classe_prevista_distancia_s1_address;       // mm_interconnect_0:PI_KNN_CLASSE_PREVISTA_DISTANCIA_s1_address -> PI_KNN_CLASSE_PREVISTA_DISTANCIA:address
	wire         mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_chipselect; // mm_interconnect_0:VGA_BUFFER_0_avalon_char_control_slave_chipselect -> VGA_BUFFER_0:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_readdata;   // VGA_BUFFER_0:ctrl_readdata -> mm_interconnect_0:VGA_BUFFER_0_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_address;    // mm_interconnect_0:VGA_BUFFER_0_avalon_char_control_slave_address -> VGA_BUFFER_0:ctrl_address
	wire         mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_read;       // mm_interconnect_0:VGA_BUFFER_0_avalon_char_control_slave_read -> VGA_BUFFER_0:ctrl_read
	wire   [3:0] mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_byteenable; // mm_interconnect_0:VGA_BUFFER_0_avalon_char_control_slave_byteenable -> VGA_BUFFER_0:ctrl_byteenable
	wire         mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_write;      // mm_interconnect_0:VGA_BUFFER_0_avalon_char_control_slave_write -> VGA_BUFFER_0:ctrl_write
	wire  [31:0] mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_writedata;  // mm_interconnect_0:VGA_BUFFER_0_avalon_char_control_slave_writedata -> VGA_BUFFER_0:ctrl_writedata
	wire         mm_interconnect_0_mmu_0_s2_chipselect;                               // mm_interconnect_0:MMU_0_s2_chipselect -> MMU_0:chipselect2
	wire  [31:0] mm_interconnect_0_mmu_0_s2_readdata;                                 // MMU_0:readdata2 -> mm_interconnect_0:MMU_0_s2_readdata
	wire   [7:0] mm_interconnect_0_mmu_0_s2_address;                                  // mm_interconnect_0:MMU_0_s2_address -> MMU_0:address2
	wire   [3:0] mm_interconnect_0_mmu_0_s2_byteenable;                               // mm_interconnect_0:MMU_0_s2_byteenable -> MMU_0:byteenable2
	wire         mm_interconnect_0_mmu_0_s2_write;                                    // mm_interconnect_0:MMU_0_s2_write -> MMU_0:write2
	wire  [31:0] mm_interconnect_0_mmu_0_s2_writedata;                                // mm_interconnect_0:MMU_0_s2_writedata -> MMU_0:writedata2
	wire         mm_interconnect_0_mmu_0_s2_clken;                                    // mm_interconnect_0:MMU_0_s2_clken -> MMU_0:clken2
	wire         irq_mapper_receiver0_irq;                                            // RS232_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                            // USB_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                            // JTAG_0:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                            // TIMER_1:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                            // TIMER_0:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_0_irq_irq;                                                     // irq_mapper:sender_irq -> NIOS2_0:irq
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [JTAG_0:rst_n, MMU_0:reset, NIOS2_0:reset_n, PIO_0:reset_n, PI_KNN_CLASSE_PREVISTA:reset_n, PI_KNN_CLASSE_PREVISTA_DISTANCIA:reset_n, PI_KNN_CLASSE_PREVISTA_PRONTO:reset_n, PO_KNN_DADOS:reset_n, PO_KNN_DADOS_ATRIBUTO:reset_n, PO_KNN_DADOS_PRONTO:reset_n, PO_KNN_K:reset_n, PO_KNN_RESET:reset_n, PO_KNN_TREINAMENTO:reset_n, RS232_0:reset, SDRAM_0:reset_n, TIMER_0:reset_n, TIMER_1:reset_n, USB_0:reset, VGA_PLL_0:reset, irq_mapper:reset, mm_interconnect_0:NIOS2_0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [MMU_0:reset_req, NIOS2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_0_debug_reset_request_reset;                                   // NIOS2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [VGA_0:reset, VGA_BUFFER_0:reset, mm_interconnect_0:VGA_BUFFER_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                  // rst_controller_002:reset_out -> [video_dual_clock_buffer_0:reset_stream_in, video_dual_clock_buffer_0:reset_stream_out]

	nios2_sopc_JTAG_0 jtag_0 (
		.clk            (clk50_0_clk),                                            //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                //               irq.irq
	);

	nios2_sopc_MMU_0 mmu_0 (
		.address     (mm_interconnect_0_mmu_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_mmu_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_mmu_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_mmu_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_mmu_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_mmu_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_mmu_0_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_mmu_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_mmu_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_mmu_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_mmu_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_mmu_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_mmu_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_mmu_0_s2_byteenable), //       .byteenable
		.clk         (clk50_0_clk),                           //   clk1.clk
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                   // (terminated)
	);

	nios2_sopc_NIOS2_0 nios2_0 (
		.clk                                 (clk50_0_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (nios2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	nios2_sopc_PIO_0 pio_0 (
		.clk        (clk50_0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)       // external_connection.export
	);

	nios2_sopc_PI_KNN_CLASSE_PREVISTA pi_knn_classe_prevista (
		.clk      (clk50_0_clk),                                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_pi_knn_classe_prevista_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pi_knn_classe_prevista_s1_readdata), //                    .readdata
		.in_port  (knn_classe_prevista_in_export)                         // external_connection.export
	);

	nios2_sopc_PI_KNN_CLASSE_PREVISTA pi_knn_classe_prevista_distancia (
		.clk      (clk50_0_clk),                                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                //               reset.reset_n
		.address  (mm_interconnect_0_pi_knn_classe_prevista_distancia_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pi_knn_classe_prevista_distancia_s1_readdata), //                    .readdata
		.in_port  (knn_classe_prevista_distancia_in_export)                         // external_connection.export
	);

	nios2_sopc_PI_KNN_CLASSE_PREVISTA_PRONTO pi_knn_classe_prevista_pronto (
		.clk      (clk50_0_clk),                                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //               reset.reset_n
		.address  (mm_interconnect_0_pi_knn_classe_prevista_pronto_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pi_knn_classe_prevista_pronto_s1_readdata), //                    .readdata
		.in_port  (knn_classe_prevista_pronto_in_export)                         // external_connection.export
	);

	nios2_sopc_PO_KNN_DADOS po_knn_dados (
		.clk        (clk50_0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_po_knn_dados_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_knn_dados_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_knn_dados_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_knn_dados_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_knn_dados_s1_readdata),   //                    .readdata
		.out_port   (knn_dados_valor_out_export)                    // external_connection.export
	);

	nios2_sopc_PO_KNN_DADOS_ATRIBUTO po_knn_dados_atributo (
		.clk        (clk50_0_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_0_po_knn_dados_atributo_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_knn_dados_atributo_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_knn_dados_atributo_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_knn_dados_atributo_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_knn_dados_atributo_s1_readdata),   //                    .readdata
		.out_port   (knn_dados_atributo_out_export)                          // external_connection.export
	);

	nios2_sopc_PO_KNN_DADOS_PRONTO po_knn_dados_pronto (
		.clk        (clk50_0_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_po_knn_dados_pronto_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_knn_dados_pronto_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_knn_dados_pronto_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_knn_dados_pronto_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_knn_dados_pronto_s1_readdata),   //                    .readdata
		.out_port   (knn_dados_pronto_out_export)                          // external_connection.export
	);

	nios2_sopc_PO_KNN_K po_knn_k (
		.clk        (clk50_0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_po_knn_k_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_knn_k_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_knn_k_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_knn_k_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_knn_k_s1_readdata),   //                    .readdata
		.out_port   (knn_k_out_export)                          // external_connection.export
	);

	nios2_sopc_PO_KNN_DADOS_PRONTO po_knn_reset (
		.clk        (clk50_0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_po_knn_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_knn_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_knn_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_knn_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_knn_reset_s1_readdata),   //                    .readdata
		.out_port   (knn_reset_out_export)                          // external_connection.export
	);

	nios2_sopc_PO_KNN_DADOS_PRONTO po_knn_treinamento (
		.clk        (clk50_0_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_po_knn_treinamento_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_knn_treinamento_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_knn_treinamento_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_knn_treinamento_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_knn_treinamento_s1_readdata),   //                    .readdata
		.out_port   (knn_treinamento_out_export)                          // external_connection.export
	);

	nios2_sopc_RS232_0 rs232_0 (
		.clk        (clk50_0_clk),                                             //                clk.clk
		.reset      (rst_controller_reset_out_reset),                          //              reset.reset
		.address    (mm_interconnect_0_rs232_0_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_rs232_0_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_rs232_0_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver0_irq),                                //          interrupt.irq
		.UART_RXD   (rs232_0_external_interface_RXD),                          // external_interface.export
		.UART_TXD   (rs232_0_external_interface_TXD)                           //                   .export
	);

	nios2_sopc_SDRAM_0 sdram_0 (
		.clk            (clk50_0_clk),                                //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),            // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                          //  wire.export
		.zs_ba          (sdram_0_wire_ba),                            //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                         //      .export
		.zs_cke         (sdram_0_wire_cke),                           //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                          //      .export
		.zs_dq          (sdram_0_wire_dq),                            //      .export
		.zs_dqm         (sdram_0_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_0_wire_we_n)                           //      .export
	);

	nios2_sopc_TIMER_0 timer_0 (
		.clk        (clk50_0_clk),                             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                 //   irq.irq
	);

	nios2_sopc_TIMER_0 timer_1 (
		.clk        (clk50_0_clk),                             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	nios2_sopc_USB_0 usb_0 (
		.clk        (clk50_0_clk),                                         //                clk.clk
		.reset      (rst_controller_reset_out_reset),                      //              reset.reset
		.address    (mm_interconnect_0_usb_0_avalon_usb_slave_address),    //   avalon_usb_slave.address
		.chipselect (mm_interconnect_0_usb_0_avalon_usb_slave_chipselect), //                   .chipselect
		.read       (mm_interconnect_0_usb_0_avalon_usb_slave_read),       //                   .read
		.write      (mm_interconnect_0_usb_0_avalon_usb_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_usb_0_avalon_usb_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_usb_0_avalon_usb_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver1_irq),                            //          interrupt.irq
		.OTG_INT1   (usb_0_external_interface_INT1),                       // external_interface.export
		.OTG_DATA   (usb_0_external_interface_DATA),                       //                   .export
		.OTG_RST_N  (usb_0_external_interface_RST_N),                      //                   .export
		.OTG_ADDR   (usb_0_external_interface_ADDR),                       //                   .export
		.OTG_CS_N   (usb_0_external_interface_CS_N),                       //                   .export
		.OTG_RD_N   (usb_0_external_interface_RD_N),                       //                   .export
		.OTG_WR_N   (usb_0_external_interface_WR_N),                       //                   .export
		.OTG_INT0   (usb_0_external_interface_INT0)                        //                   .export
	);

	nios2_sopc_VGA_0 vga_0 (
		.clk           (vga_pll_0_c0_clk),                                                //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                              //              reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_0_external_interface_CLK),                                    // external_interface.export
		.VGA_HS        (vga_0_external_interface_HS),                                     //                   .export
		.VGA_VS        (vga_0_external_interface_VS),                                     //                   .export
		.VGA_BLANK     (vga_0_external_interface_BLANK),                                  //                   .export
		.VGA_SYNC      (vga_0_external_interface_SYNC),                                   //                   .export
		.VGA_R         (vga_0_external_interface_R),                                      //                   .export
		.VGA_G         (vga_0_external_interface_G),                                      //                   .export
		.VGA_B         (vga_0_external_interface_B)                                       //                   .export
	);

	nios2_sopc_VGA_BUFFER_0 vga_buffer_0 (
		.clk                  (vga_pll_0_c0_clk),                                                    //                       clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                  //                     reset.reset
		.ctrl_address         (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (vga_buffer_0_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (vga_buffer_0_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (vga_buffer_0_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (vga_buffer_0_avalon_char_source_valid),                               //                          .valid
		.stream_data          (vga_buffer_0_avalon_char_source_data)                                 //                          .data
	);

	nios2_sopc_VGA_PLL_0 vga_pll_0 (
		.clk                (clk50_0_clk),                                     //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read               (mm_interconnect_0_vga_pll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_vga_pll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_vga_pll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_vga_pll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_vga_pll_0_pll_slave_writedata), //                      .writedata
		.c0                 (vga_pll_0_c0_clk),                                //                    c0.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (4'b0000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	nios2_sopc_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (vga_pll_0_c0_clk),                                                //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_002_reset_out_reset),                              //         reset_stream_in.reset
		.clk_stream_out           (vga_pll_0_c0_clk),                                                //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                              //        reset_stream_out.reset
		.stream_in_ready          (vga_buffer_0_avalon_char_source_ready),                           //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (vga_buffer_0_avalon_char_source_startofpacket),                   //                        .startofpacket
		.stream_in_endofpacket    (vga_buffer_0_avalon_char_source_endofpacket),                     //                        .endofpacket
		.stream_in_valid          (vga_buffer_0_avalon_char_source_valid),                           //                        .valid
		.stream_in_data           (vga_buffer_0_avalon_char_source_data),                            //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	nios2_sopc_mm_interconnect_0 mm_interconnect_0 (
		.CLK50_0_clk_clk                                   (clk50_0_clk),                                                         //                              CLK50_0_clk.clk
		.VGA_PLL_0_c0_clk                                  (vga_pll_0_c0_clk),                                                    //                             VGA_PLL_0_c0.clk
		.NIOS2_0_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                      //      NIOS2_0_reset_reset_bridge_in_reset.reset
		.VGA_BUFFER_0_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                                  // VGA_BUFFER_0_reset_reset_bridge_in_reset.reset
		.NIOS2_0_data_master_address                       (nios2_0_data_master_address),                                         //                      NIOS2_0_data_master.address
		.NIOS2_0_data_master_waitrequest                   (nios2_0_data_master_waitrequest),                                     //                                         .waitrequest
		.NIOS2_0_data_master_byteenable                    (nios2_0_data_master_byteenable),                                      //                                         .byteenable
		.NIOS2_0_data_master_read                          (nios2_0_data_master_read),                                            //                                         .read
		.NIOS2_0_data_master_readdata                      (nios2_0_data_master_readdata),                                        //                                         .readdata
		.NIOS2_0_data_master_readdatavalid                 (nios2_0_data_master_readdatavalid),                                   //                                         .readdatavalid
		.NIOS2_0_data_master_write                         (nios2_0_data_master_write),                                           //                                         .write
		.NIOS2_0_data_master_writedata                     (nios2_0_data_master_writedata),                                       //                                         .writedata
		.NIOS2_0_data_master_debugaccess                   (nios2_0_data_master_debugaccess),                                     //                                         .debugaccess
		.NIOS2_0_instruction_master_address                (nios2_0_instruction_master_address),                                  //               NIOS2_0_instruction_master.address
		.NIOS2_0_instruction_master_waitrequest            (nios2_0_instruction_master_waitrequest),                              //                                         .waitrequest
		.NIOS2_0_instruction_master_read                   (nios2_0_instruction_master_read),                                     //                                         .read
		.NIOS2_0_instruction_master_readdata               (nios2_0_instruction_master_readdata),                                 //                                         .readdata
		.NIOS2_0_instruction_master_readdatavalid          (nios2_0_instruction_master_readdatavalid),                            //                                         .readdatavalid
		.JTAG_0_avalon_jtag_slave_address                  (mm_interconnect_0_jtag_0_avalon_jtag_slave_address),                  //                 JTAG_0_avalon_jtag_slave.address
		.JTAG_0_avalon_jtag_slave_write                    (mm_interconnect_0_jtag_0_avalon_jtag_slave_write),                    //                                         .write
		.JTAG_0_avalon_jtag_slave_read                     (mm_interconnect_0_jtag_0_avalon_jtag_slave_read),                     //                                         .read
		.JTAG_0_avalon_jtag_slave_readdata                 (mm_interconnect_0_jtag_0_avalon_jtag_slave_readdata),                 //                                         .readdata
		.JTAG_0_avalon_jtag_slave_writedata                (mm_interconnect_0_jtag_0_avalon_jtag_slave_writedata),                //                                         .writedata
		.JTAG_0_avalon_jtag_slave_waitrequest              (mm_interconnect_0_jtag_0_avalon_jtag_slave_waitrequest),              //                                         .waitrequest
		.JTAG_0_avalon_jtag_slave_chipselect               (mm_interconnect_0_jtag_0_avalon_jtag_slave_chipselect),               //                                         .chipselect
		.MMU_0_s1_address                                  (mm_interconnect_0_mmu_0_s1_address),                                  //                                 MMU_0_s1.address
		.MMU_0_s1_write                                    (mm_interconnect_0_mmu_0_s1_write),                                    //                                         .write
		.MMU_0_s1_readdata                                 (mm_interconnect_0_mmu_0_s1_readdata),                                 //                                         .readdata
		.MMU_0_s1_writedata                                (mm_interconnect_0_mmu_0_s1_writedata),                                //                                         .writedata
		.MMU_0_s1_byteenable                               (mm_interconnect_0_mmu_0_s1_byteenable),                               //                                         .byteenable
		.MMU_0_s1_chipselect                               (mm_interconnect_0_mmu_0_s1_chipselect),                               //                                         .chipselect
		.MMU_0_s1_clken                                    (mm_interconnect_0_mmu_0_s1_clken),                                    //                                         .clken
		.MMU_0_s2_address                                  (mm_interconnect_0_mmu_0_s2_address),                                  //                                 MMU_0_s2.address
		.MMU_0_s2_write                                    (mm_interconnect_0_mmu_0_s2_write),                                    //                                         .write
		.MMU_0_s2_readdata                                 (mm_interconnect_0_mmu_0_s2_readdata),                                 //                                         .readdata
		.MMU_0_s2_writedata                                (mm_interconnect_0_mmu_0_s2_writedata),                                //                                         .writedata
		.MMU_0_s2_byteenable                               (mm_interconnect_0_mmu_0_s2_byteenable),                               //                                         .byteenable
		.MMU_0_s2_chipselect                               (mm_interconnect_0_mmu_0_s2_chipselect),                               //                                         .chipselect
		.MMU_0_s2_clken                                    (mm_interconnect_0_mmu_0_s2_clken),                                    //                                         .clken
		.NIOS2_0_debug_mem_slave_address                   (mm_interconnect_0_nios2_0_debug_mem_slave_address),                   //                  NIOS2_0_debug_mem_slave.address
		.NIOS2_0_debug_mem_slave_write                     (mm_interconnect_0_nios2_0_debug_mem_slave_write),                     //                                         .write
		.NIOS2_0_debug_mem_slave_read                      (mm_interconnect_0_nios2_0_debug_mem_slave_read),                      //                                         .read
		.NIOS2_0_debug_mem_slave_readdata                  (mm_interconnect_0_nios2_0_debug_mem_slave_readdata),                  //                                         .readdata
		.NIOS2_0_debug_mem_slave_writedata                 (mm_interconnect_0_nios2_0_debug_mem_slave_writedata),                 //                                         .writedata
		.NIOS2_0_debug_mem_slave_byteenable                (mm_interconnect_0_nios2_0_debug_mem_slave_byteenable),                //                                         .byteenable
		.NIOS2_0_debug_mem_slave_waitrequest               (mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest),               //                                         .waitrequest
		.NIOS2_0_debug_mem_slave_debugaccess               (mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess),               //                                         .debugaccess
		.PI_KNN_CLASSE_PREVISTA_s1_address                 (mm_interconnect_0_pi_knn_classe_prevista_s1_address),                 //                PI_KNN_CLASSE_PREVISTA_s1.address
		.PI_KNN_CLASSE_PREVISTA_s1_readdata                (mm_interconnect_0_pi_knn_classe_prevista_s1_readdata),                //                                         .readdata
		.PI_KNN_CLASSE_PREVISTA_DISTANCIA_s1_address       (mm_interconnect_0_pi_knn_classe_prevista_distancia_s1_address),       //      PI_KNN_CLASSE_PREVISTA_DISTANCIA_s1.address
		.PI_KNN_CLASSE_PREVISTA_DISTANCIA_s1_readdata      (mm_interconnect_0_pi_knn_classe_prevista_distancia_s1_readdata),      //                                         .readdata
		.PI_KNN_CLASSE_PREVISTA_PRONTO_s1_address          (mm_interconnect_0_pi_knn_classe_prevista_pronto_s1_address),          //         PI_KNN_CLASSE_PREVISTA_PRONTO_s1.address
		.PI_KNN_CLASSE_PREVISTA_PRONTO_s1_readdata         (mm_interconnect_0_pi_knn_classe_prevista_pronto_s1_readdata),         //                                         .readdata
		.PIO_0_s1_address                                  (mm_interconnect_0_pio_0_s1_address),                                  //                                 PIO_0_s1.address
		.PIO_0_s1_write                                    (mm_interconnect_0_pio_0_s1_write),                                    //                                         .write
		.PIO_0_s1_readdata                                 (mm_interconnect_0_pio_0_s1_readdata),                                 //                                         .readdata
		.PIO_0_s1_writedata                                (mm_interconnect_0_pio_0_s1_writedata),                                //                                         .writedata
		.PIO_0_s1_chipselect                               (mm_interconnect_0_pio_0_s1_chipselect),                               //                                         .chipselect
		.PO_KNN_DADOS_s1_address                           (mm_interconnect_0_po_knn_dados_s1_address),                           //                          PO_KNN_DADOS_s1.address
		.PO_KNN_DADOS_s1_write                             (mm_interconnect_0_po_knn_dados_s1_write),                             //                                         .write
		.PO_KNN_DADOS_s1_readdata                          (mm_interconnect_0_po_knn_dados_s1_readdata),                          //                                         .readdata
		.PO_KNN_DADOS_s1_writedata                         (mm_interconnect_0_po_knn_dados_s1_writedata),                         //                                         .writedata
		.PO_KNN_DADOS_s1_chipselect                        (mm_interconnect_0_po_knn_dados_s1_chipselect),                        //                                         .chipselect
		.PO_KNN_DADOS_ATRIBUTO_s1_address                  (mm_interconnect_0_po_knn_dados_atributo_s1_address),                  //                 PO_KNN_DADOS_ATRIBUTO_s1.address
		.PO_KNN_DADOS_ATRIBUTO_s1_write                    (mm_interconnect_0_po_knn_dados_atributo_s1_write),                    //                                         .write
		.PO_KNN_DADOS_ATRIBUTO_s1_readdata                 (mm_interconnect_0_po_knn_dados_atributo_s1_readdata),                 //                                         .readdata
		.PO_KNN_DADOS_ATRIBUTO_s1_writedata                (mm_interconnect_0_po_knn_dados_atributo_s1_writedata),                //                                         .writedata
		.PO_KNN_DADOS_ATRIBUTO_s1_chipselect               (mm_interconnect_0_po_knn_dados_atributo_s1_chipselect),               //                                         .chipselect
		.PO_KNN_DADOS_PRONTO_s1_address                    (mm_interconnect_0_po_knn_dados_pronto_s1_address),                    //                   PO_KNN_DADOS_PRONTO_s1.address
		.PO_KNN_DADOS_PRONTO_s1_write                      (mm_interconnect_0_po_knn_dados_pronto_s1_write),                      //                                         .write
		.PO_KNN_DADOS_PRONTO_s1_readdata                   (mm_interconnect_0_po_knn_dados_pronto_s1_readdata),                   //                                         .readdata
		.PO_KNN_DADOS_PRONTO_s1_writedata                  (mm_interconnect_0_po_knn_dados_pronto_s1_writedata),                  //                                         .writedata
		.PO_KNN_DADOS_PRONTO_s1_chipselect                 (mm_interconnect_0_po_knn_dados_pronto_s1_chipselect),                 //                                         .chipselect
		.PO_KNN_K_s1_address                               (mm_interconnect_0_po_knn_k_s1_address),                               //                              PO_KNN_K_s1.address
		.PO_KNN_K_s1_write                                 (mm_interconnect_0_po_knn_k_s1_write),                                 //                                         .write
		.PO_KNN_K_s1_readdata                              (mm_interconnect_0_po_knn_k_s1_readdata),                              //                                         .readdata
		.PO_KNN_K_s1_writedata                             (mm_interconnect_0_po_knn_k_s1_writedata),                             //                                         .writedata
		.PO_KNN_K_s1_chipselect                            (mm_interconnect_0_po_knn_k_s1_chipselect),                            //                                         .chipselect
		.PO_KNN_RESET_s1_address                           (mm_interconnect_0_po_knn_reset_s1_address),                           //                          PO_KNN_RESET_s1.address
		.PO_KNN_RESET_s1_write                             (mm_interconnect_0_po_knn_reset_s1_write),                             //                                         .write
		.PO_KNN_RESET_s1_readdata                          (mm_interconnect_0_po_knn_reset_s1_readdata),                          //                                         .readdata
		.PO_KNN_RESET_s1_writedata                         (mm_interconnect_0_po_knn_reset_s1_writedata),                         //                                         .writedata
		.PO_KNN_RESET_s1_chipselect                        (mm_interconnect_0_po_knn_reset_s1_chipselect),                        //                                         .chipselect
		.PO_KNN_TREINAMENTO_s1_address                     (mm_interconnect_0_po_knn_treinamento_s1_address),                     //                    PO_KNN_TREINAMENTO_s1.address
		.PO_KNN_TREINAMENTO_s1_write                       (mm_interconnect_0_po_knn_treinamento_s1_write),                       //                                         .write
		.PO_KNN_TREINAMENTO_s1_readdata                    (mm_interconnect_0_po_knn_treinamento_s1_readdata),                    //                                         .readdata
		.PO_KNN_TREINAMENTO_s1_writedata                   (mm_interconnect_0_po_knn_treinamento_s1_writedata),                   //                                         .writedata
		.PO_KNN_TREINAMENTO_s1_chipselect                  (mm_interconnect_0_po_knn_treinamento_s1_chipselect),                  //                                         .chipselect
		.RS232_0_avalon_rs232_slave_address                (mm_interconnect_0_rs232_0_avalon_rs232_slave_address),                //               RS232_0_avalon_rs232_slave.address
		.RS232_0_avalon_rs232_slave_write                  (mm_interconnect_0_rs232_0_avalon_rs232_slave_write),                  //                                         .write
		.RS232_0_avalon_rs232_slave_read                   (mm_interconnect_0_rs232_0_avalon_rs232_slave_read),                   //                                         .read
		.RS232_0_avalon_rs232_slave_readdata               (mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata),               //                                         .readdata
		.RS232_0_avalon_rs232_slave_writedata              (mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata),              //                                         .writedata
		.RS232_0_avalon_rs232_slave_byteenable             (mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable),             //                                         .byteenable
		.RS232_0_avalon_rs232_slave_chipselect             (mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect),             //                                         .chipselect
		.SDRAM_0_s1_address                                (mm_interconnect_0_sdram_0_s1_address),                                //                               SDRAM_0_s1.address
		.SDRAM_0_s1_write                                  (mm_interconnect_0_sdram_0_s1_write),                                  //                                         .write
		.SDRAM_0_s1_read                                   (mm_interconnect_0_sdram_0_s1_read),                                   //                                         .read
		.SDRAM_0_s1_readdata                               (mm_interconnect_0_sdram_0_s1_readdata),                               //                                         .readdata
		.SDRAM_0_s1_writedata                              (mm_interconnect_0_sdram_0_s1_writedata),                              //                                         .writedata
		.SDRAM_0_s1_byteenable                             (mm_interconnect_0_sdram_0_s1_byteenable),                             //                                         .byteenable
		.SDRAM_0_s1_readdatavalid                          (mm_interconnect_0_sdram_0_s1_readdatavalid),                          //                                         .readdatavalid
		.SDRAM_0_s1_waitrequest                            (mm_interconnect_0_sdram_0_s1_waitrequest),                            //                                         .waitrequest
		.SDRAM_0_s1_chipselect                             (mm_interconnect_0_sdram_0_s1_chipselect),                             //                                         .chipselect
		.TIMER_0_s1_address                                (mm_interconnect_0_timer_0_s1_address),                                //                               TIMER_0_s1.address
		.TIMER_0_s1_write                                  (mm_interconnect_0_timer_0_s1_write),                                  //                                         .write
		.TIMER_0_s1_readdata                               (mm_interconnect_0_timer_0_s1_readdata),                               //                                         .readdata
		.TIMER_0_s1_writedata                              (mm_interconnect_0_timer_0_s1_writedata),                              //                                         .writedata
		.TIMER_0_s1_chipselect                             (mm_interconnect_0_timer_0_s1_chipselect),                             //                                         .chipselect
		.TIMER_1_s1_address                                (mm_interconnect_0_timer_1_s1_address),                                //                               TIMER_1_s1.address
		.TIMER_1_s1_write                                  (mm_interconnect_0_timer_1_s1_write),                                  //                                         .write
		.TIMER_1_s1_readdata                               (mm_interconnect_0_timer_1_s1_readdata),                               //                                         .readdata
		.TIMER_1_s1_writedata                              (mm_interconnect_0_timer_1_s1_writedata),                              //                                         .writedata
		.TIMER_1_s1_chipselect                             (mm_interconnect_0_timer_1_s1_chipselect),                             //                                         .chipselect
		.USB_0_avalon_usb_slave_address                    (mm_interconnect_0_usb_0_avalon_usb_slave_address),                    //                   USB_0_avalon_usb_slave.address
		.USB_0_avalon_usb_slave_write                      (mm_interconnect_0_usb_0_avalon_usb_slave_write),                      //                                         .write
		.USB_0_avalon_usb_slave_read                       (mm_interconnect_0_usb_0_avalon_usb_slave_read),                       //                                         .read
		.USB_0_avalon_usb_slave_readdata                   (mm_interconnect_0_usb_0_avalon_usb_slave_readdata),                   //                                         .readdata
		.USB_0_avalon_usb_slave_writedata                  (mm_interconnect_0_usb_0_avalon_usb_slave_writedata),                  //                                         .writedata
		.USB_0_avalon_usb_slave_chipselect                 (mm_interconnect_0_usb_0_avalon_usb_slave_chipselect),                 //                                         .chipselect
		.VGA_BUFFER_0_avalon_char_buffer_slave_address     (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_address),     //    VGA_BUFFER_0_avalon_char_buffer_slave.address
		.VGA_BUFFER_0_avalon_char_buffer_slave_write       (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_write),       //                                         .write
		.VGA_BUFFER_0_avalon_char_buffer_slave_read        (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_read),        //                                         .read
		.VGA_BUFFER_0_avalon_char_buffer_slave_readdata    (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_readdata),    //                                         .readdata
		.VGA_BUFFER_0_avalon_char_buffer_slave_writedata   (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_writedata),   //                                         .writedata
		.VGA_BUFFER_0_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_byteenable),  //                                         .byteenable
		.VGA_BUFFER_0_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_waitrequest), //                                         .waitrequest
		.VGA_BUFFER_0_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_vga_buffer_0_avalon_char_buffer_slave_chipselect),  //                                         .chipselect
		.VGA_BUFFER_0_avalon_char_control_slave_address    (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_address),    //   VGA_BUFFER_0_avalon_char_control_slave.address
		.VGA_BUFFER_0_avalon_char_control_slave_write      (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_write),      //                                         .write
		.VGA_BUFFER_0_avalon_char_control_slave_read       (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_read),       //                                         .read
		.VGA_BUFFER_0_avalon_char_control_slave_readdata   (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_readdata),   //                                         .readdata
		.VGA_BUFFER_0_avalon_char_control_slave_writedata  (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_writedata),  //                                         .writedata
		.VGA_BUFFER_0_avalon_char_control_slave_byteenable (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_byteenable), //                                         .byteenable
		.VGA_BUFFER_0_avalon_char_control_slave_chipselect (mm_interconnect_0_vga_buffer_0_avalon_char_control_slave_chipselect), //                                         .chipselect
		.VGA_PLL_0_pll_slave_address                       (mm_interconnect_0_vga_pll_0_pll_slave_address),                       //                      VGA_PLL_0_pll_slave.address
		.VGA_PLL_0_pll_slave_write                         (mm_interconnect_0_vga_pll_0_pll_slave_write),                         //                                         .write
		.VGA_PLL_0_pll_slave_read                          (mm_interconnect_0_vga_pll_0_pll_slave_read),                          //                                         .read
		.VGA_PLL_0_pll_slave_readdata                      (mm_interconnect_0_vga_pll_0_pll_slave_readdata),                      //                                         .readdata
		.VGA_PLL_0_pll_slave_writedata                     (mm_interconnect_0_vga_pll_0_pll_slave_writedata)                      //                                         .writedata
	);

	nios2_sopc_irq_mapper irq_mapper (
		.clk           (clk50_0_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_0_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_clk50_0_reset_n),             // reset_in0.reset
		.reset_in1      (nios2_0_debug_reset_request_reset),  // reset_in1.reset
		.clk            (clk50_0_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_clk50_0_reset_n),             // reset_in0.reset
		.reset_in1      (nios2_0_debug_reset_request_reset),  // reset_in1.reset
		.clk            (vga_pll_0_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_clk50_0_reset_n),             // reset_in0.reset
		.clk            (vga_pll_0_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
