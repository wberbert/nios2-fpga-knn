library ieee;
use ieee.std_logic_1164.all;

package berbert_parallel_buble_sort_type is

end package berbert_parallel_buble_sort_type;

library ieee;
use ieee.std_logic_1164.all;
use work.lcd_types.all;