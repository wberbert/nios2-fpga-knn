-- nios2_sopc.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios2_sopc is
	port (
		clk50_0_clk                      : in    std_logic                     := '0';             --                    clk50_0.clk
		pio_0_external_connection_export : out   std_logic_vector(7 downto 0);                     --  pio_0_external_connection.export
		reset_clk50_0_reset_n            : in    std_logic                     := '0';             --              reset_clk50_0.reset_n
		rs232_0_external_interface_RXD   : in    std_logic                     := '0';             -- rs232_0_external_interface.RXD
		rs232_0_external_interface_TXD   : out   std_logic;                                        --                           .TXD
		sdram_0_wire_addr                : out   std_logic_vector(12 downto 0);                    --               sdram_0_wire.addr
		sdram_0_wire_ba                  : out   std_logic_vector(1 downto 0);                     --                           .ba
		sdram_0_wire_cas_n               : out   std_logic;                                        --                           .cas_n
		sdram_0_wire_cke                 : out   std_logic;                                        --                           .cke
		sdram_0_wire_cs_n                : out   std_logic;                                        --                           .cs_n
		sdram_0_wire_dq                  : inout std_logic_vector(31 downto 0) := (others => '0'); --                           .dq
		sdram_0_wire_dqm                 : out   std_logic_vector(3 downto 0);                     --                           .dqm
		sdram_0_wire_ras_n               : out   std_logic;                                        --                           .ras_n
		sdram_0_wire_we_n                : out   std_logic                                         --                           .we_n
	);
end entity nios2_sopc;

architecture rtl of nios2_sopc is
	component nios2_sopc_JTAG_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios2_sopc_JTAG_0;

	component nios2_sopc_MMU_0 is
		port (
			address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component nios2_sopc_MMU_0;

	component nios2_sopc_NIOS2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios2_sopc_NIOS2_0;

	component nios2_sopc_PIO_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios2_sopc_PIO_0;

	component nios2_sopc_RS232_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic                     := 'X';             -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			irq        : out std_logic;                                        -- irq
			UART_RXD   : in  std_logic                     := 'X';             -- export
			UART_TXD   : out std_logic                                         -- export
		);
	end component nios2_sopc_RS232_0;

	component nios2_sopc_SDRAM_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios2_sopc_SDRAM_0;

	component nios2_sopc_TIMER_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios2_sopc_TIMER_0;

	component nios2_sopc_mm_interconnect_0 is
		port (
			CLK50_0_clk_clk                           : in  std_logic                     := 'X';             -- clk
			NIOS2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			NIOS2_0_data_master_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			NIOS2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			NIOS2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOS2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			NIOS2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS2_0_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			NIOS2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			NIOS2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOS2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			NIOS2_0_instruction_master_address        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			NIOS2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			NIOS2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			NIOS2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS2_0_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			JTAG_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			JTAG_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			JTAG_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			JTAG_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			JTAG_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			MMU_0_s1_address                          : out std_logic_vector(7 downto 0);                     -- address
			MMU_0_s1_write                            : out std_logic;                                        -- write
			MMU_0_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			MMU_0_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			MMU_0_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			MMU_0_s1_chipselect                       : out std_logic;                                        -- chipselect
			MMU_0_s1_clken                            : out std_logic;                                        -- clken
			MMU_0_s2_address                          : out std_logic_vector(7 downto 0);                     -- address
			MMU_0_s2_write                            : out std_logic;                                        -- write
			MMU_0_s2_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			MMU_0_s2_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			MMU_0_s2_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			MMU_0_s2_chipselect                       : out std_logic;                                        -- chipselect
			MMU_0_s2_clken                            : out std_logic;                                        -- clken
			NIOS2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			NIOS2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			NIOS2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			NIOS2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOS2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			NIOS2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOS2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			NIOS2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			PIO_0_s1_address                          : out std_logic_vector(2 downto 0);                     -- address
			PIO_0_s1_write                            : out std_logic;                                        -- write
			PIO_0_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PIO_0_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			PIO_0_s1_chipselect                       : out std_logic;                                        -- chipselect
			RS232_0_avalon_rs232_slave_address        : out std_logic_vector(0 downto 0);                     -- address
			RS232_0_avalon_rs232_slave_write          : out std_logic;                                        -- write
			RS232_0_avalon_rs232_slave_read           : out std_logic;                                        -- read
			RS232_0_avalon_rs232_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RS232_0_avalon_rs232_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			RS232_0_avalon_rs232_slave_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			RS232_0_avalon_rs232_slave_chipselect     : out std_logic;                                        -- chipselect
			SDRAM_0_s1_address                        : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_0_s1_write                          : out std_logic;                                        -- write
			SDRAM_0_s1_read                           : out std_logic;                                        -- read
			SDRAM_0_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SDRAM_0_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			SDRAM_0_s1_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			SDRAM_0_s1_readdatavalid                  : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_0_s1_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_0_s1_chipselect                     : out std_logic;                                        -- chipselect
			TIMER_0_s1_address                        : out std_logic_vector(2 downto 0);                     -- address
			TIMER_0_s1_write                          : out std_logic;                                        -- write
			TIMER_0_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			TIMER_0_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			TIMER_0_s1_chipselect                     : out std_logic;                                        -- chipselect
			TIMER_1_s1_address                        : out std_logic_vector(2 downto 0);                     -- address
			TIMER_1_s1_write                          : out std_logic;                                        -- write
			TIMER_1_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			TIMER_1_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			TIMER_1_s1_chipselect                     : out std_logic                                         -- chipselect
		);
	end component nios2_sopc_mm_interconnect_0;

	component nios2_sopc_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios2_sopc_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_0_data_master_readdata -> NIOS2_0:d_readdata
	signal nios2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:NIOS2_0_data_master_waitrequest -> NIOS2_0:d_waitrequest
	signal nios2_0_data_master_debugaccess                            : std_logic;                     -- NIOS2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_0_data_master_debugaccess
	signal nios2_0_data_master_address                                : std_logic_vector(27 downto 0); -- NIOS2_0:d_address -> mm_interconnect_0:NIOS2_0_data_master_address
	signal nios2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- NIOS2_0:d_byteenable -> mm_interconnect_0:NIOS2_0_data_master_byteenable
	signal nios2_0_data_master_read                                   : std_logic;                     -- NIOS2_0:d_read -> mm_interconnect_0:NIOS2_0_data_master_read
	signal nios2_0_data_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:NIOS2_0_data_master_readdatavalid -> NIOS2_0:d_readdatavalid
	signal nios2_0_data_master_write                                  : std_logic;                     -- NIOS2_0:d_write -> mm_interconnect_0:NIOS2_0_data_master_write
	signal nios2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- NIOS2_0:d_writedata -> mm_interconnect_0:NIOS2_0_data_master_writedata
	signal nios2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_0_instruction_master_readdata -> NIOS2_0:i_readdata
	signal nios2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:NIOS2_0_instruction_master_waitrequest -> NIOS2_0:i_waitrequest
	signal nios2_0_instruction_master_address                         : std_logic_vector(27 downto 0); -- NIOS2_0:i_address -> mm_interconnect_0:NIOS2_0_instruction_master_address
	signal nios2_0_instruction_master_read                            : std_logic;                     -- NIOS2_0:i_read -> mm_interconnect_0:NIOS2_0_instruction_master_read
	signal nios2_0_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:NIOS2_0_instruction_master_readdatavalid -> NIOS2_0:i_readdatavalid
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_0_avalon_jtag_slave_chipselect -> JTAG_0:av_chipselect
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_0:av_readdata -> mm_interconnect_0:JTAG_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_0:av_waitrequest -> mm_interconnect_0:JTAG_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_0_avalon_jtag_slave_address -> JTAG_0:av_address
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_0_avalon_jtag_slave_writedata -> JTAG_0:av_writedata
	signal mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect    : std_logic;                     -- mm_interconnect_0:RS232_0_avalon_rs232_slave_chipselect -> RS232_0:chipselect
	signal mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata      : std_logic_vector(31 downto 0); -- RS232_0:readdata -> mm_interconnect_0:RS232_0_avalon_rs232_slave_readdata
	signal mm_interconnect_0_rs232_0_avalon_rs232_slave_address       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:RS232_0_avalon_rs232_slave_address -> RS232_0:address
	signal mm_interconnect_0_rs232_0_avalon_rs232_slave_read          : std_logic;                     -- mm_interconnect_0:RS232_0_avalon_rs232_slave_read -> RS232_0:read
	signal mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RS232_0_avalon_rs232_slave_byteenable -> RS232_0:byteenable
	signal mm_interconnect_0_rs232_0_avalon_rs232_slave_write         : std_logic;                     -- mm_interconnect_0:RS232_0_avalon_rs232_slave_write -> RS232_0:write
	signal mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:RS232_0_avalon_rs232_slave_writedata -> RS232_0:writedata
	signal mm_interconnect_0_nios2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- NIOS2_0:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest      : std_logic;                     -- NIOS2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:NIOS2_0_debug_mem_slave_debugaccess -> NIOS2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NIOS2_0_debug_mem_slave_address -> NIOS2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:NIOS2_0_debug_mem_slave_read -> NIOS2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NIOS2_0_debug_mem_slave_byteenable -> NIOS2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:NIOS2_0_debug_mem_slave_write -> NIOS2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_0_debug_mem_slave_writedata -> NIOS2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_mmu_0_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:MMU_0_s1_chipselect -> MMU_0:chipselect
	signal mm_interconnect_0_mmu_0_s1_readdata                        : std_logic_vector(31 downto 0); -- MMU_0:readdata -> mm_interconnect_0:MMU_0_s1_readdata
	signal mm_interconnect_0_mmu_0_s1_address                         : std_logic_vector(7 downto 0);  -- mm_interconnect_0:MMU_0_s1_address -> MMU_0:address
	signal mm_interconnect_0_mmu_0_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:MMU_0_s1_byteenable -> MMU_0:byteenable
	signal mm_interconnect_0_mmu_0_s1_write                           : std_logic;                     -- mm_interconnect_0:MMU_0_s1_write -> MMU_0:write
	signal mm_interconnect_0_mmu_0_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:MMU_0_s1_writedata -> MMU_0:writedata
	signal mm_interconnect_0_mmu_0_s1_clken                           : std_logic;                     -- mm_interconnect_0:MMU_0_s1_clken -> MMU_0:clken
	signal mm_interconnect_0_sdram_0_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:SDRAM_0_s1_chipselect -> SDRAM_0:az_cs
	signal mm_interconnect_0_sdram_0_s1_readdata                      : std_logic_vector(31 downto 0); -- SDRAM_0:za_data -> mm_interconnect_0:SDRAM_0_s1_readdata
	signal mm_interconnect_0_sdram_0_s1_waitrequest                   : std_logic;                     -- SDRAM_0:za_waitrequest -> mm_interconnect_0:SDRAM_0_s1_waitrequest
	signal mm_interconnect_0_sdram_0_s1_address                       : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_0_s1_address -> SDRAM_0:az_addr
	signal mm_interconnect_0_sdram_0_s1_read                          : std_logic;                     -- mm_interconnect_0:SDRAM_0_s1_read -> mm_interconnect_0_sdram_0_s1_read:in
	signal mm_interconnect_0_sdram_0_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SDRAM_0_s1_byteenable -> mm_interconnect_0_sdram_0_s1_byteenable:in
	signal mm_interconnect_0_sdram_0_s1_readdatavalid                 : std_logic;                     -- SDRAM_0:za_valid -> mm_interconnect_0:SDRAM_0_s1_readdatavalid
	signal mm_interconnect_0_sdram_0_s1_write                         : std_logic;                     -- mm_interconnect_0:SDRAM_0_s1_write -> mm_interconnect_0_sdram_0_s1_write:in
	signal mm_interconnect_0_sdram_0_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:SDRAM_0_s1_writedata -> SDRAM_0:az_data
	signal mm_interconnect_0_pio_0_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:PIO_0_s1_chipselect -> PIO_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                        : std_logic_vector(31 downto 0); -- PIO_0:readdata -> mm_interconnect_0:PIO_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:PIO_0_s1_address -> PIO_0:address
	signal mm_interconnect_0_pio_0_s1_write                           : std_logic;                     -- mm_interconnect_0:PIO_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:PIO_0_s1_writedata -> PIO_0:writedata
	signal mm_interconnect_0_timer_1_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:TIMER_1_s1_chipselect -> TIMER_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                      : std_logic_vector(15 downto 0); -- TIMER_1:readdata -> mm_interconnect_0:TIMER_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TIMER_1_s1_address -> TIMER_1:address
	signal mm_interconnect_0_timer_1_s1_write                         : std_logic;                     -- mm_interconnect_0:TIMER_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:TIMER_1_s1_writedata -> TIMER_1:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:TIMER_0_s1_chipselect -> TIMER_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                      : std_logic_vector(15 downto 0); -- TIMER_0:readdata -> mm_interconnect_0:TIMER_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TIMER_0_s1_address -> TIMER_0:address
	signal mm_interconnect_0_timer_0_s1_write                         : std_logic;                     -- mm_interconnect_0:TIMER_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:TIMER_0_s1_writedata -> TIMER_0:writedata
	signal mm_interconnect_0_mmu_0_s2_chipselect                      : std_logic;                     -- mm_interconnect_0:MMU_0_s2_chipselect -> MMU_0:chipselect2
	signal mm_interconnect_0_mmu_0_s2_readdata                        : std_logic_vector(31 downto 0); -- MMU_0:readdata2 -> mm_interconnect_0:MMU_0_s2_readdata
	signal mm_interconnect_0_mmu_0_s2_address                         : std_logic_vector(7 downto 0);  -- mm_interconnect_0:MMU_0_s2_address -> MMU_0:address2
	signal mm_interconnect_0_mmu_0_s2_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:MMU_0_s2_byteenable -> MMU_0:byteenable2
	signal mm_interconnect_0_mmu_0_s2_write                           : std_logic;                     -- mm_interconnect_0:MMU_0_s2_write -> MMU_0:write2
	signal mm_interconnect_0_mmu_0_s2_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:MMU_0_s2_writedata -> MMU_0:writedata2
	signal mm_interconnect_0_mmu_0_s2_clken                           : std_logic;                     -- mm_interconnect_0:MMU_0_s2_clken -> MMU_0:clken2
	signal irq_mapper_receiver0_irq                                   : std_logic;                     -- RS232_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                   : std_logic;                     -- JTAG_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                   : std_logic;                     -- TIMER_1:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                   : std_logic;                     -- TIMER_0:irq -> irq_mapper:receiver3_irq
	signal nios2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NIOS2_0:irq
	signal rst_controller_reset_out_reset                             : std_logic;                     -- rst_controller:reset_out -> [MMU_0:reset, RS232_0:reset, irq_mapper:reset, mm_interconnect_0:NIOS2_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                         : std_logic;                     -- rst_controller:reset_req -> [MMU_0:reset_req, NIOS2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_0_debug_reset_request_reset                          : std_logic;                     -- NIOS2_0:debug_reset_request -> rst_controller:reset_in1
	signal reset_clk50_0_reset_n_ports_inv                            : std_logic;                     -- reset_clk50_0_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_0_avalon_jtag_slave_read:inv -> JTAG_0:av_read_n
	signal mm_interconnect_0_jtag_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_0_avalon_jtag_slave_write:inv -> JTAG_0:av_write_n
	signal mm_interconnect_0_sdram_0_s1_read_ports_inv                : std_logic;                     -- mm_interconnect_0_sdram_0_s1_read:inv -> SDRAM_0:az_rd_n
	signal mm_interconnect_0_sdram_0_s1_byteenable_ports_inv          : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_0_s1_byteenable:inv -> SDRAM_0:az_be_n
	signal mm_interconnect_0_sdram_0_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_sdram_0_s1_write:inv -> SDRAM_0:az_wr_n
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> PIO_0:write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> TIMER_1:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> TIMER_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JTAG_0:rst_n, NIOS2_0:reset_n, PIO_0:reset_n, SDRAM_0:reset_n, TIMER_0:reset_n, TIMER_1:reset_n]

begin

	jtag_0 : component nios2_sopc_JTAG_0
		port map (
			clk            => clk50_0_clk,                                                --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                   --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                    --               irq.irq
		);

	mmu_0 : component nios2_sopc_MMU_0
		port map (
			address     => mm_interconnect_0_mmu_0_s1_address,    --     s1.address
			clken       => mm_interconnect_0_mmu_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_mmu_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_mmu_0_s1_write,      --       .write
			readdata    => mm_interconnect_0_mmu_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_mmu_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_mmu_0_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_0_mmu_0_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_mmu_0_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_mmu_0_s2_clken,      --       .clken
			write2      => mm_interconnect_0_mmu_0_s2_write,      --       .write
			readdata2   => mm_interconnect_0_mmu_0_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_mmu_0_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_mmu_0_s2_byteenable, --       .byteenable
			clk         => clk50_0_clk,                           --   clk1.clk
			reset       => rst_controller_reset_out_reset,        -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,    --       .reset_req
			freeze      => '0'                                    -- (terminated)
		);

	nios2_0 : component nios2_sopc_NIOS2_0
		port map (
			clk                                 => clk50_0_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,              --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                           => nios2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	pio_0 : component nios2_sopc_PIO_0
		port map (
			clk        => clk50_0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			out_port   => pio_0_external_connection_export            -- external_connection.export
		);

	rs232_0 : component nios2_sopc_RS232_0
		port map (
			clk        => clk50_0_clk,                                             --                clk.clk
			reset      => rst_controller_reset_out_reset,                          --              reset.reset
			address    => mm_interconnect_0_rs232_0_avalon_rs232_slave_address(0), -- avalon_rs232_slave.address
			chipselect => mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect, --                   .chipselect
			byteenable => mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable, --                   .byteenable
			read       => mm_interconnect_0_rs232_0_avalon_rs232_slave_read,       --                   .read
			write      => mm_interconnect_0_rs232_0_avalon_rs232_slave_write,      --                   .write
			writedata  => mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata,  --                   .writedata
			readdata   => mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata,   --                   .readdata
			irq        => irq_mapper_receiver0_irq,                                --          interrupt.irq
			UART_RXD   => rs232_0_external_interface_RXD,                          -- external_interface.export
			UART_TXD   => rs232_0_external_interface_TXD                           --                   .export
		);

	sdram_0 : component nios2_sopc_SDRAM_0
		port map (
			clk            => clk50_0_clk,                                       --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,          -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_0_wire_addr,                                 --  wire.export
			zs_ba          => sdram_0_wire_ba,                                   --      .export
			zs_cas_n       => sdram_0_wire_cas_n,                                --      .export
			zs_cke         => sdram_0_wire_cke,                                  --      .export
			zs_cs_n        => sdram_0_wire_cs_n,                                 --      .export
			zs_dq          => sdram_0_wire_dq,                                   --      .export
			zs_dqm         => sdram_0_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_0_wire_ras_n,                                --      .export
			zs_we_n        => sdram_0_wire_we_n                                  --      .export
		);

	timer_0 : component nios2_sopc_TIMER_0
		port map (
			clk        => clk50_0_clk,                                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                      --   irq.irq
		);

	timer_1 : component nios2_sopc_TIMER_0
		port map (
			clk        => clk50_0_clk,                                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                      --   irq.irq
		);

	mm_interconnect_0 : component nios2_sopc_mm_interconnect_0
		port map (
			CLK50_0_clk_clk                           => clk50_0_clk,                                             --                         CLK50_0_clk.clk
			NIOS2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                          -- NIOS2_0_reset_reset_bridge_in_reset.reset
			NIOS2_0_data_master_address               => nios2_0_data_master_address,                             --                 NIOS2_0_data_master.address
			NIOS2_0_data_master_waitrequest           => nios2_0_data_master_waitrequest,                         --                                    .waitrequest
			NIOS2_0_data_master_byteenable            => nios2_0_data_master_byteenable,                          --                                    .byteenable
			NIOS2_0_data_master_read                  => nios2_0_data_master_read,                                --                                    .read
			NIOS2_0_data_master_readdata              => nios2_0_data_master_readdata,                            --                                    .readdata
			NIOS2_0_data_master_readdatavalid         => nios2_0_data_master_readdatavalid,                       --                                    .readdatavalid
			NIOS2_0_data_master_write                 => nios2_0_data_master_write,                               --                                    .write
			NIOS2_0_data_master_writedata             => nios2_0_data_master_writedata,                           --                                    .writedata
			NIOS2_0_data_master_debugaccess           => nios2_0_data_master_debugaccess,                         --                                    .debugaccess
			NIOS2_0_instruction_master_address        => nios2_0_instruction_master_address,                      --          NIOS2_0_instruction_master.address
			NIOS2_0_instruction_master_waitrequest    => nios2_0_instruction_master_waitrequest,                  --                                    .waitrequest
			NIOS2_0_instruction_master_read           => nios2_0_instruction_master_read,                         --                                    .read
			NIOS2_0_instruction_master_readdata       => nios2_0_instruction_master_readdata,                     --                                    .readdata
			NIOS2_0_instruction_master_readdatavalid  => nios2_0_instruction_master_readdatavalid,                --                                    .readdatavalid
			JTAG_0_avalon_jtag_slave_address          => mm_interconnect_0_jtag_0_avalon_jtag_slave_address,      --            JTAG_0_avalon_jtag_slave.address
			JTAG_0_avalon_jtag_slave_write            => mm_interconnect_0_jtag_0_avalon_jtag_slave_write,        --                                    .write
			JTAG_0_avalon_jtag_slave_read             => mm_interconnect_0_jtag_0_avalon_jtag_slave_read,         --                                    .read
			JTAG_0_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_0_avalon_jtag_slave_readdata,     --                                    .readdata
			JTAG_0_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_0_avalon_jtag_slave_writedata,    --                                    .writedata
			JTAG_0_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_0_avalon_jtag_slave_waitrequest,  --                                    .waitrequest
			JTAG_0_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_0_avalon_jtag_slave_chipselect,   --                                    .chipselect
			MMU_0_s1_address                          => mm_interconnect_0_mmu_0_s1_address,                      --                            MMU_0_s1.address
			MMU_0_s1_write                            => mm_interconnect_0_mmu_0_s1_write,                        --                                    .write
			MMU_0_s1_readdata                         => mm_interconnect_0_mmu_0_s1_readdata,                     --                                    .readdata
			MMU_0_s1_writedata                        => mm_interconnect_0_mmu_0_s1_writedata,                    --                                    .writedata
			MMU_0_s1_byteenable                       => mm_interconnect_0_mmu_0_s1_byteenable,                   --                                    .byteenable
			MMU_0_s1_chipselect                       => mm_interconnect_0_mmu_0_s1_chipselect,                   --                                    .chipselect
			MMU_0_s1_clken                            => mm_interconnect_0_mmu_0_s1_clken,                        --                                    .clken
			MMU_0_s2_address                          => mm_interconnect_0_mmu_0_s2_address,                      --                            MMU_0_s2.address
			MMU_0_s2_write                            => mm_interconnect_0_mmu_0_s2_write,                        --                                    .write
			MMU_0_s2_readdata                         => mm_interconnect_0_mmu_0_s2_readdata,                     --                                    .readdata
			MMU_0_s2_writedata                        => mm_interconnect_0_mmu_0_s2_writedata,                    --                                    .writedata
			MMU_0_s2_byteenable                       => mm_interconnect_0_mmu_0_s2_byteenable,                   --                                    .byteenable
			MMU_0_s2_chipselect                       => mm_interconnect_0_mmu_0_s2_chipselect,                   --                                    .chipselect
			MMU_0_s2_clken                            => mm_interconnect_0_mmu_0_s2_clken,                        --                                    .clken
			NIOS2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_0_debug_mem_slave_address,       --             NIOS2_0_debug_mem_slave.address
			NIOS2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_0_debug_mem_slave_write,         --                                    .write
			NIOS2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_0_debug_mem_slave_read,          --                                    .read
			NIOS2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_0_debug_mem_slave_readdata,      --                                    .readdata
			NIOS2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_0_debug_mem_slave_writedata,     --                                    .writedata
			NIOS2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_0_debug_mem_slave_byteenable,    --                                    .byteenable
			NIOS2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest,   --                                    .waitrequest
			NIOS2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess,   --                                    .debugaccess
			PIO_0_s1_address                          => mm_interconnect_0_pio_0_s1_address,                      --                            PIO_0_s1.address
			PIO_0_s1_write                            => mm_interconnect_0_pio_0_s1_write,                        --                                    .write
			PIO_0_s1_readdata                         => mm_interconnect_0_pio_0_s1_readdata,                     --                                    .readdata
			PIO_0_s1_writedata                        => mm_interconnect_0_pio_0_s1_writedata,                    --                                    .writedata
			PIO_0_s1_chipselect                       => mm_interconnect_0_pio_0_s1_chipselect,                   --                                    .chipselect
			RS232_0_avalon_rs232_slave_address        => mm_interconnect_0_rs232_0_avalon_rs232_slave_address,    --          RS232_0_avalon_rs232_slave.address
			RS232_0_avalon_rs232_slave_write          => mm_interconnect_0_rs232_0_avalon_rs232_slave_write,      --                                    .write
			RS232_0_avalon_rs232_slave_read           => mm_interconnect_0_rs232_0_avalon_rs232_slave_read,       --                                    .read
			RS232_0_avalon_rs232_slave_readdata       => mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata,   --                                    .readdata
			RS232_0_avalon_rs232_slave_writedata      => mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata,  --                                    .writedata
			RS232_0_avalon_rs232_slave_byteenable     => mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable, --                                    .byteenable
			RS232_0_avalon_rs232_slave_chipselect     => mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect, --                                    .chipselect
			SDRAM_0_s1_address                        => mm_interconnect_0_sdram_0_s1_address,                    --                          SDRAM_0_s1.address
			SDRAM_0_s1_write                          => mm_interconnect_0_sdram_0_s1_write,                      --                                    .write
			SDRAM_0_s1_read                           => mm_interconnect_0_sdram_0_s1_read,                       --                                    .read
			SDRAM_0_s1_readdata                       => mm_interconnect_0_sdram_0_s1_readdata,                   --                                    .readdata
			SDRAM_0_s1_writedata                      => mm_interconnect_0_sdram_0_s1_writedata,                  --                                    .writedata
			SDRAM_0_s1_byteenable                     => mm_interconnect_0_sdram_0_s1_byteenable,                 --                                    .byteenable
			SDRAM_0_s1_readdatavalid                  => mm_interconnect_0_sdram_0_s1_readdatavalid,              --                                    .readdatavalid
			SDRAM_0_s1_waitrequest                    => mm_interconnect_0_sdram_0_s1_waitrequest,                --                                    .waitrequest
			SDRAM_0_s1_chipselect                     => mm_interconnect_0_sdram_0_s1_chipselect,                 --                                    .chipselect
			TIMER_0_s1_address                        => mm_interconnect_0_timer_0_s1_address,                    --                          TIMER_0_s1.address
			TIMER_0_s1_write                          => mm_interconnect_0_timer_0_s1_write,                      --                                    .write
			TIMER_0_s1_readdata                       => mm_interconnect_0_timer_0_s1_readdata,                   --                                    .readdata
			TIMER_0_s1_writedata                      => mm_interconnect_0_timer_0_s1_writedata,                  --                                    .writedata
			TIMER_0_s1_chipselect                     => mm_interconnect_0_timer_0_s1_chipselect,                 --                                    .chipselect
			TIMER_1_s1_address                        => mm_interconnect_0_timer_1_s1_address,                    --                          TIMER_1_s1.address
			TIMER_1_s1_write                          => mm_interconnect_0_timer_1_s1_write,                      --                                    .write
			TIMER_1_s1_readdata                       => mm_interconnect_0_timer_1_s1_readdata,                   --                                    .readdata
			TIMER_1_s1_writedata                      => mm_interconnect_0_timer_1_s1_writedata,                  --                                    .writedata
			TIMER_1_s1_chipselect                     => mm_interconnect_0_timer_1_s1_chipselect                  --                                    .chipselect
		);

	irq_mapper : component nios2_sopc_irq_mapper
		port map (
			clk           => clk50_0_clk,                    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_0_irq_irq                 --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_clk50_0_reset_n_ports_inv,    -- reset_in0.reset
			reset_in1      => nios2_0_debug_reset_request_reset,  -- reset_in1.reset
			clk            => clk50_0_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_clk50_0_reset_n_ports_inv <= not reset_clk50_0_reset_n;

	mm_interconnect_0_jtag_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_0_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_0_s1_read_ports_inv <= not mm_interconnect_0_sdram_0_s1_read;

	mm_interconnect_0_sdram_0_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_0_s1_byteenable;

	mm_interconnect_0_sdram_0_s1_write_ports_inv <= not mm_interconnect_0_sdram_0_s1_write;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios2_sopc
